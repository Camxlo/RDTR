library verilog;
use verilog.vl_types.all;
entity Mod6 is
    port(
        Q0              : out    vl_logic;
        Entrada         : in     vl_logic;
        Q1              : out    vl_logic;
        Q2              : out    vl_logic
    );
end Mod6;
