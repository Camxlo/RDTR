library verilog;
use verilog.vl_types.all;
entity Mod6_vlg_vec_tst is
end Mod6_vlg_vec_tst;
