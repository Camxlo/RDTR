library verilog;
use verilog.vl_types.all;
entity Mod6_vlg_sample_tst is
    port(
        Entrada         : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Mod6_vlg_sample_tst;
